module hazard_unit(
      input wire [31:0] instruction_ID_EX,
      input wire [4:0] rd_EX_MEM,
      input wire mem_read_ID_EX,
      output reg pc_write,
      output reg IF_ID_write
   );


always @(*) begin
   
end
   
endmodule

